library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity full_adder IS
port (
      a,b,cin :in std_logic_vector(0 downto 0);
      sum,carry : out STD_LOGIC
      );
end entity;

architecture behavioral of full_adder is

signal s1 : std_logic_vector(1 downto 0);

begin
      process (a,b,cin)
      begin
        s1 <= ('0'& a) + ('0'& b) +('0'& cin);
      
      end process;
      carry <= s1(1);
      sum <= s1(0);

end architecture;
