library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;


entity ask2 is 

    generic (
        
    );
    port (

    );

end entity;


architecture behavioral of ask2 is 
    signal 

    begin 

    process (clock,reset)

    end process;

    
end architecture;